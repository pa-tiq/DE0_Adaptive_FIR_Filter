LIBRARY work;
USE work.constants_and_types.ALL;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fir_filter_lms_test is
	generic( 
		BUTTON_HIGH 	: STD_LOGIC := '0' );
	port (
		clk              	  : in  std_logic;
		reset                 : in  std_logic;
		o_data_buffer         : out OUT_TYPE;
		o_fir_coeff1          : out IN_TYPE;
		o_fir_coeff2          : out IN_TYPE;
		o_inputref		      : out IN_TYPE;
		o_inputdata		      : out IN_TYPE;
		o_error               : out OUT_TYPE);
end fir_filter_lms_test;

architecture rtl of fir_filter_lms_test is

	--x = [64,111,-64,-111,64,111,-64,-111,64,111,-64,-111,64,111,-64];
	--d = [10,60,9,-41,10,60,10,-39,11,60,10,-40,10,59,9];
	--y = [-7,-1,5,20,-9,-36,5,40,-8,-50,2,48,-4,-53,-1,49,-3,-52];
	
	constant noisy_size : integer := 15;
	type T_NOISY_INPUT is array(0 to noisy_size-1) of integer range (-2**Win) to (2**Win-1);
	type T_COEFF_INPUT is array(0 to LFilter-1) of integer range (-2**Win) to (2**Win-1);

	constant NOISY_ARRAY : T_NOISY_INPUT := (
		64,111,-64,-111,64,111,-64,-111,64,111,-64,-111,64,111,-64
	);
	constant NOISYF_ARRAY : T_NOISY_INPUT := (
		10,60,9,-41,10,60,10,-39,11,60,10,-40,10,59,9
	);

	-- degrau tamanho 512
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	0,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- degrau tamanho 1024
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	0,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,
	--	255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);

	-- noisy sin -127 to 126
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-10,1,11,35,36,18,49,41,42,51,51,56,70,75,79,79,72,87,96,93,100,
	--	101,98,104,100,111,101,103,106,95,121,115,109,121,103,111,109,111,
	--	110,101,104,101,103,103,100,85,87,76,73,75,80,62,64,56,59,41,42,40,
	--	38,35,21,6,5,-3,11,-11,-9,-20,-19,-35,-44,-49,-43,-52,-58,-53,-64,
	--	-70,-66,-84,-80,-83,-93,-93,-105,-108,-103,-102,-94,-114,-111,-114,
	--	-126,-119,-127,-112,-122,-117,-120,-114);

	--noisy sawtooth -64 to 63
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-30,-25,-33,-32,-20,-46,-30,-35,-26,-15,-12,-27,-20,-13,-15,-8 ,-6 ,-16,-8 ,-24,7  ,-7 ,-11,0  ,-9 ,5  ,2  ,28 ,20 ,-11,17 ,2  ,14 ,19 ,26 ,19 ,37 ,20 ,29 ,33 ,30 ,39 ,35 ,27 ,19 ,54 ,33 ,41 ,47 ,44 ,37 ,42 ,47 ,63 ,44 ,60 ,57 ,54 ,48 ,57 ,60 ,50 ,-35,-42,-34,-29,-38,-31,-24,-42,-14,0  ,-12,-22,-13,-25,3  ,-4 ,-4 ,-17,-5 ,-11,-7 ,-8 ,-10,-8 ,0  ,-12,11 ,6  ,15 ,13 ,16 ,0  ,6  ,12 ,19 ,30 ,19 ,34
	--	);

	--noisy sawtooth -256 to 255
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	-155,-124,-155,-177,-200,-134,-104,-138,-140,-125,-147,-119,-102,-87 ,-85 ,-54 ,-65 ,2   ,-45 ,15  ,-70 ,-18 ,-40 ,-3  ,3   ,-90 ,-53 ,-50 ,22  ,67  ,9   ,56  ,53  ,2   ,61  ,26  ,114 ,64  ,131 ,63  ,106 ,89  ,25  ,69  ,133 ,115 ,83  ,107 ,145 ,107 ,184 ,132 ,227 ,130 ,182 ,127 ,162 ,173 ,215 ,241 ,224 ,206 ,256 ,-142,-160,-138,-137,-181,-112,-156,-148,-113,-124,-112,-79 ,-56 ,-95 ,-69 ,-83 ,-60 ,-46 ,-78 ,-39 ,-21 ,-33 ,32  ,-45 ,-43 ,-73 ,29  ,34  ,6   ,48  ,28  ,39  ,39  ,57  ,51  ,154 ,18		
	--);

	-- TAMANHO 1060 - Símbolo OFDM parte real, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,-8,-252,-50,257,131,-90,5,157,127,28,-93,-149,13,112,-163,-382,-122,189,158,75,50,-166,-386,-280,-62,56,178,156,-138,-239,35,83,-201,-143,231,201,-134,-148,1,-117,-248,-126,-9,2,87,129,-59,-271,-297,-202,-33,141,83,-163,-215,-66,-97,-263,-163,123,159,-20,-31,131,200,217,341,368,100,-137,-28,131,38,-18,179,270,60,-114,-110,-115,-81,52,-8,-247,-187,132,176,39,121,92,-338,-512,-44,336,189,63,176,112,-90,-67,20,-13,69,172,-87,-376,-133,229,58,-304,-288,-133,-161,-152,-17,-24,-148,-149,-103,-160,-203,-158,-129,-90,43,175,221,202,51,-220,-289,-14,210,91,-72,3,85,-48,-167,-25,196,187,-7,-75,77,226,197,58,-77,-135,-26,191,227,19,-99,13,48,-119,-185,-14,138,105,-7,-104,-172,-151,2,184,210,29,-159,-169,-116,-120,-8,225,186,-104,-43,339,272,-225,-285,114,187,-14,158,477,337,16,45,179,45,-156,-171,-75,31,77,-34,-202,-229,-164,-112,-2,112,34,-119,-49,160,181,4,-106,-8,186,250,115,-8,-1,-61,-202,-102,179,155,-121,-81,239,290,115,159,267,41,-228,-63,287,284,-20,-204,-157,-101,-174,-232,-56,255,328,94,-53,36,11,-217,-228,49,140,-45,-60,109,12,-313,-394,-226,-153,-178,-138,-96,-73,16,11,-215,-365,-244,-130,-145,-76,-21,-204,-296,-6,207,-5,-209,-135,-115,-189,-86,-34,-244,-209,268,447,71,-90,178,183,-131,-134,82,-16,-223,-157,-133,-348,-375,-130,-45,-77,99,201,-86,-292,-7,338,313,117,-46,-220,-281,-96,99,58,-109,-215,-183,-6,125,-24,-241,-108,242,305,42,-131,-13,202,265,149,52,97,127,35,-9,56,57,36,179,300,140,-77,-95,-73,-87,46,211,125,-25,51,150,39,-51,65,170,68,-127,-204,-96,53,96,145,303,322,100,17,194,195,-36,-18,230,190,-114,-226,-86,105,261,236,-21,-195,-152,-181,-259,-17,368,361,41,-120,-67,-9,-6,-78,-192,-174,-20,54,55,143,232,174,56,-12,-31,-25,-94,-263,-259,57,301,220,109,115,43,-34,58,80,-61,3,278,314,123,46,8,-77,3,84,-165,-312,105,468,163,-240,-149,16,-107,-151,49,138,24,-13,76,92,-11,-104,-147,-217,-276,-153,82,98,-75,-58,66,-105,-355,-225,-21,-172,-298,-93,-26,-247,-185,209,309,60,-46,9,-52,-124,-38,49,49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- TAMANHO 1060 - Símbolo OFDM parte imaginária, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,-241,-142,-79,-110,-46,-71,-296,-384,-232,-109,17,300,443,217,-3,66,131,-16,-132,-64,31,78,150,181,59,-55,59,201,8,-327,-267,80,90,-225,-240,70,115,-147,-184,64,136,-73,-201,-68,116,121,0,-46,19,12,-155,-341,-401,-342,-250,-197,-172,-110,-78,-175,-203,51,280,108,-189,-172,11,80,137,199,80,-51,88,265,191,87,129,79,-124,-203,-104,-26,-33,-85,-129,-47,129,164,58,44,92,53,53,139,59,-177,-251,-176,-158,-81,88,14,-268,-254,66,195,108,138,211,138,91,111,-100,-466,-465,-32,262,78,-250,-268,-3,153,26,-161,-198,-138,-45,63,35,-146,-126,222,407,129,-168,-117,-36,-211,-380,-298,-89,106,239,191,-11,-91,29,102,24,-58,-112,-179,-112,128,206,-49,-245,-59,190,133,-14,73,212,114,-108,-231,-248,-160,38,128,-31,-134,26,87,-180,-350,-147,-1,-217,-432,-339,-134,-5,125,246,217,47,-112,-151,-115,-150,-249,-210,-77,-146,-270,1,405,262,-189,-178,118,30,-220,-79,180,106,-79,-106,-112,-141,-93,-51,-13,198,425,308,-20,-125,29,162,122,-38,-135,-34,128,186,215,202,4,-107,199,465,137,-321,-258,49,127,67,-36,-198,-147,139,143,-155,-187,-4,-83,-227,-121,-98,-266,-193,34,-35,-163,6,139,66,144,279,76,-185,-129,-73,-194,-162,-40,-181,-347,-180,102,270,382,335,142,165,312,96,-219,-43,238,11,-296,-145,99,97,97,106,-101,-281,-154,1,-66,-142,-47,142,258,89,-318,-436,-27,333,196,-58,-33,86,98,61,-7,-83,-31,102,105,-3,-60,-55,-31,-10,-72,-175,-106,94,120,-28,-69,-15,-49,-51,124,265,197,122,168,114,-152,-357,-266,-73,-69,-142,35,376,419,67,-220,-125,122,213,154,76,51,108,171,117,12,36,128,87,-17,32,175,182,32,-132,-231,-230,-128,-16,67,138,56,-250,-368,3,302,-23,-363,13,511,294,-139,22,371,226,-92,-65,70,9,-45,59,143,127,98,97,136,167,34,-227,-286,-46,137,26,-140,-81,110,140,-56,-232,-165,50,170,133,23,-87,-110,-14,66,45,69,205,223,-28,-320,-322,2,349,374,100,-83,5,79,-58,-176,-73,124,234,216,98,-15,-33,-59,-171,-187,-22,53,-71,-95,90,156,-9,-79,48,69,-82,-88,92,94,-162,-316,-222,-113,-105,-108,-92,-7,200,271,-5,-199,70,278,-47,-332,-62,265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- A saída da convolução vai ter tamanho 1572

	-- TAMANHO 1060 - Símbolo OFDM parte real, -1024 to 1023
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	97,213,470,554,368,99,-75,-138,-167,-126,10,-63,-548,-931,-650,-34,246,143,34,99,196,68,-202,-139,221,205,-161,-76,428,620,556,552,211,-348,-240,237,-17,-504,-99,513,263,-180,10,314,253,56,-186,-298,26,225,-325,-764,-243,378,316,150,100,-333,-771,-561,-123,113,356,311,-275,-478,69,166,-403,-285,463,402,-269,-295,2,-234,-497,-251,-17,3,174,258,-118,-543,-594,-404,-65,282,166,-326,-430,-131,-194,-527,-326,246,318,-41,-63,262,400,434,682,735,201,-274,-56,263,76,-36,358,539,120,-228,-220,-230,-162,103,-15,-495,-373,265,352,78,242,185,-676,-1024,-88,671,379,126,352,224,-179,-135,40,-27,138,344,-174,-751,-266,458,115,-607,-576,-266,-323,-303,-34,-47,-295,-299,-207,-321,-405,-315,-257,-180,85,350,442,404,102,-439,-578,-28,421,183,-144,5,170,-96,-333,-50,392,373,-13,-150,154,452,394,115,-153,-271,-51,383,455,38,-198,25,96,-237,-370,-29,276,210,-14,-207,-343,-302,3,368,419,59,-317,-339,-232,-241,-16,450,371,-208,-86,678,543,-451,-571,228,374,-28,316,955,673,32,90,359,90,-313,-343,-151,62,154,-68,-403,-458,-328,-224,-4,224,68,-238,-97,320,362,9,-211,-16,373,500,229,-15,-1,-121,-403,-204,358,309,-241,-162,479,581,230,319,534,83,-456,-125,574,569,-39,-408,-315,-202,-348,-464,-112,511,655,188,-107,72,22,-434,-457,99,279,-91,-121,219,23,-627,-789,-451,-306,-356,-275,-193,-146,32,22,-431,-731,-487,-260,-290,-152,-43,-409,-593,-13,414,-10,-418,-271,-231,-378,-173,-68,-489,-418,536,894,142,-181,356,366,-262,-268,164,-33,-446,-314,-266,-697,-750,-260,-90,-154,199,402,-172,-584,-14,676,627,233,-92,-440,-563,-192,197,116,-219,-430,-366,-13,250,-48,-482,-216,483,609,83,-262,-25,405,530,298,105,194,254,71,-18,112,114,73,359,599,280,-155,-190,-146,-174,93,421,250,-50,103,299,77,-102,131,340,136,-254,-408,-193,105,191,291,605,645,201,34,388,390,-73,-36,459,380,-227,-452,-172,211,523,472,-42,-391,-305,-362,-518,-34,736,722,82,-240,-133,-19,-13,-155,-384,-347,-40,109,110,285,464,349,111,-24,-61,-50,-187,-527,-517,115,602,441,217,231,87,-67,115,160,-123,6,557,628,247,92,16,-154,6,167,-329,-623,210,936,325,-480,-299,32,-213,-302,98,275,47,-26,152,184,-21,-207,-293,-433,-552,-305,165,197,-150,-117,133,-210,-709,-450,-42,-343,-595,-186,-52,-495,-370,419,619,120,-92,19,-105,-248,-76,97,97,213,470,554,368,99,-75,-138,-167,-126,10,-63,-548,-931,-650,-34,246,143,34,99,196,68,-202,-139,221,205,-161,-76,428,620,556,552,211,-348,-240,237,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- TAMANHO 1060 - Símbolo OFDM parte imaginária, -1024 to 1023
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	530,470,334,262,-238,-476,236,783,330,-60,175,119,-249,17,584,518,136,4,-97,-103,275,438,-82,-500,-239,111,103,-27,-101,-3,282,221,-319,-358,399,681,0,-482,-285,-158,-221,-92,-142,-592,-768,-465,-218,35,601,886,434,-7,131,262,-31,-264,-128,62,155,300,362,118,-109,118,403,16,-654,-536,159,179,-450,-480,141,230,-295,-369,128,272,-146,-403,-136,231,243,0,-91,38,24,-311,-682,-802,-685,-500,-394,-344,-220,-156,-350,-406,102,561,216,-379,-344,21,159,274,398,160,-102,175,530,383,173,258,159,-248,-406,-208,-52,-67,-170,-258,-94,258,328,117,88,184,106,106,278,118,-355,-502,-352,-317,-163,177,29,-537,-508,132,391,217,276,422,276,181,222,-200,-933,-931,-63,525,156,-501,-536,-7,306,51,-322,-397,-277,-90,127,70,-293,-253,444,815,258,-337,-234,-72,-423,-761,-596,-179,212,478,381,-22,-182,59,205,48,-117,-225,-358,-224,255,412,-99,-490,-118,381,265,-27,146,425,229,-216,-463,-497,-321,77,256,-62,-268,51,174,-361,-700,-294,-2,-434,-866,-678,-269,-11,251,492,434,94,-223,-302,-230,-300,-498,-421,-155,-292,-541,3,812,525,-378,-356,236,59,-440,-158,360,213,-159,-212,-223,-283,-187,-102,-26,397,851,616,-40,-250,59,325,245,-77,-271,-68,257,372,430,404,8,-214,399,930,275,-642,-517,98,254,133,-71,-397,-293,278,286,-310,-374,-9,-166,-454,-242,-196,-533,-387,67,-71,-326,12,279,131,288,558,151,-370,-259,-145,-389,-324,-80,-361,-694,-360,205,541,765,670,284,331,626,193,-439,-86,476,21,-593,-290,197,195,194,213,-202,-563,-308,1,-132,-284,-93,284,517,177,-637,-873,-54,667,393,-115,-67,173,196,122,-13,-165,-62,203,211,-6,-121,-110,-62,-20,-143,-350,-212,188,240,-56,-139,-30,-98,-102,249,530,395,244,336,229,-305,-714,-532,-146,-138,-284,70,752,839,133,-439,-250,244,427,309,152,102,216,342,234,24,72,256,175,-33,65,350,364,65,-264,-463,-461,-257,-31,134,277,112,-500,-738,6,605,-46,-727,25,1023,588,-278,43,743,452,-184,-131,139,17,-89,118,287,254,196,195,273,335,68,-455,-573,-93,273,52,-281,-161,219,280,-112,-464,-329,99,339,266,45,-174,-220,-28,133,90,137,409,447,-56,-640,-645,3,699,748,199,-165,11,157,-116,-353,-146,248,469,433,196,-30,-66,-118,-343,-373,-44,106,-143,-191,179,312,-17,-159,96,138,-164,-175,185,188,-324,-633,-445,-226,-210,-216,-185,-14,401,543,-11,-399,139,557,-93,-665,-125,530,470,334,262,-238,-476,236,783,330,-60,175,119,-249,17,584,518,136,4,-97,-103,275,438,-82,-500,-239,111,103,-27,-101,-3,282,221,-319,-358,399,681,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- A saída da convolução vai ter tamanho 1572, mas só preciso dos 1060

	--------------------------------------------------------------------
	-- TAMANHO 1060 - Símbolo OFDM filtrado parte real, -1024 to 1023
	--constant NOISYF_ARRAY : T_NOISY_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,0,-1,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,2,-1,-1,1,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,2,-2,-1,2,-1,-2,2,1,-2,1,2,-2,-1,3,0,-2,2,1,-3,0,3,-2,-2,3,0,-3,2,2,-3,0,3,-2,-2,3,0,-3,2,2,-4,0,4,-2,-3,4,1,-4,2,3,-4,-1,5,-2,-4,5,1,-5,2,4,-5,-2,6,-2,-5,5,2,-6,1,3,6,74,244,454,545,388,92,-87,-124,-167,-139,18,-56,-559,-930,-640,-41,241,152,32,91,203,71,-210,-138,228,200,-164,-69,427,614,561,554,205,-347,-235,233,-19,-499,-100,509,266,-178,5,315,258,53,-188,-294,26,221,-323,-762,-247,379,320,148,98,-330,-771,-564,-121,115,354,311,-273,-480,67,168,-403,-288,464,404,-271,-296,5,-235,-499,-249,-17,1,175,260,-120,-544,-592,-405,-67,284,167,-329,-429,-130,-195,-528,-324,246,317,-40,-62,261,401,436,681,735,202,-274,-58,264,77,-38,358,541,120,-229,-218,-229,-163,104,-15,-496,-374,266,352,77,243,185,-677,-1024,-87,671,378,127,352,223,-179,-135,39,-26,139,344,-174,-751,-266,458,116,-607,-577,-266,-322,-304,-35,-46,-295,-299,-206,-320,-406,-315,-257,-180,85,351,442,403,102,-439,-579,-28,422,183,-145,6,171,-96,-333,-49,392,373,-13,-150,154,453,394,115,-153,-271,-51,383,455,38,-198,26,96,-238,-370,-29,276,210,-14,-207,-343,-302,3,367,419,59,-317,-339,-232,-241,-17,450,372,-208,-86,679,544,-451,-571,228,374,-28,316,955,673,32,90,359,90,-313,-343,-151,62,154,-68,-403,-458,-328,-224,-4,224,68,-238,-97,320,362,9,-211,-16,373,500,229,-15,-1,-121,-403,-204,358,310,-241,-162,479,581,230,319,534,83,-456,-125,574,569,-39,-408,-315,-202,-348,-464,-112,511,655,188,-106,72,22,-434,-457,99,280,-91,-121,219,24,-627,-789,-451,-306,-356,-275,-193,-147,32,22,-431,-731,-488,-260,-290,-152,-43,-409,-593,-13,414,-10,-418,-271,-231,-378,-173,-69,-489,-418,536,894,143,-181,356,367,-262,-269,164,-32,-446,-315,-266,-697,-751,-260,-90,-154,199,402,-173,-584,-14,676,627,233,-92,-441,-563,-192,197,115,-218,-430,-367,-12,250,-48,-482,-215,483,609,84,-262,-26,405,530,297,105,195,254,70,-17,113,113,73,360,599,280,-154,-190,-147,-174,93,420,251,-49,102,299,79,-103,130,341,137,-255,-408,-192,104,191,293,605,643,202,35,386,390,-71,-37,458,381,-227,-454,-171,212,521,471,-39,-392,-307,-361,-517,-37,737,725,80,-241,-130,-19,-15,-154,-383,-350,-40,112,108,284,467,349,108,-22,-59,-53,-187,-523,-520,113,606,441,213,233,89,-71,115,165,-125,2,561,629,243,93,20,-158,5,173,-331,-628,215,939,320,-479,-294,28,-216,-296,97,270,52,-23,146,184,-15,-212,-297,-426,-553,-312,169,202,-158,-117,141,-214,-715,-442,-42,-352,-591,-179,-60,-496,-360,414,611,129,-90,8,-100,-239,-86,94,110,208,459,566,372,84,-70,-126,-181,-131,28,-68,-563,-916,-643,-55,251,161,16,90,222,61,-226,-116,232,172,-151,-44,396,606,606,532,164,-283,-229,124,138,-62,-35,60,-9,-41,30,16,-35,6,27,-21,-12,25,-4,-20,16,10,-20,3,17,-12,-9,16,-2,-14,10,8,-14,1,13,-8,-7,12,0,-11,7,7,-10,-1,10,-5,-7,9,1,-9,4,6,-8,-1,8,-3,-6,7,2,-8,3,6,-6,-2,7,-2,-5,5,2,-6,1,5,-4,-3,6,-1,-5,4,3,-5,1,5,-3,-3,5,0,-4,3,3,-4,0,4,-2,-3,4,0,-4,2,3,-3,-1,3,-1,-3,3,1,-3,1,3,-2,-1,3,-1,-2,2,1,-3,1,2,-2,-1,2,0,-2,2,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,0,2,-1,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
	--);
	-- TAMANHO 1060 - Símbolo OFDM filtrado parte imaginária, -1024 to 1023
	--constant NOISYF_ARRAY : T_NOISY_INPUT := (
	--	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,-1,0,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,1,-2,0,1,-1,-1,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-2,0,2,-1,-2,2,0,-3,1,2,-2,0,3,-1,-2,3,1,-3,1,3,-3,-1,3,-1,-3,3,1,-4,1,3,-3,-2,4,-1,-4,3,2,-4,0,4,-3,-3,5,0,-5,3,3,-5,0,5,-3,-4,5,1,-6,3,4,-6,-1,7,-3,-5,6,2,-7,3,6,-6,-2,8,-2,-7,7,3,-9,2,8,-7,-4,10,-2,-9,8,5,-11,2,11,-8,-6,13,-1,-13,9,8,-14,1,15,-10,-9,17,-1,-18,12,12,-20,0,22,-15,-15,26,0,-29,20,20,-36,2,42,-32,-29,64,-12,-94,148,438,457,404,228,-268,-433,234,749,352,-44,147,121,-225,2,572,539,135,-14,-86,-93,259,439,-67,-509,-249,124,104,-39,-94,5,272,221,-309,-363,392,691,2,-492,-281,-152,-229,-94,-134,-596,-776,-459,-216,27,604,893,429,-9,138,261,-37,-259,-125,56,157,305,358,116,-104,117,398,20,-652,-541,160,184,-454,-483,145,231,-300,-367,131,268,-147,-399,-138,229,247,0,-95,40,27,-314,-684,-800,-688,-504,-392,-343,-223,-156,-348,-409,101,565,215,-382,-343,22,157,275,401,159,-103,178,531,381,175,260,157,-248,-405,-209,-53,-65,-170,-260,-93,260,327,117,90,184,105,107,279,116,-355,-502,-354,-318,-161,176,28,-537,-508,131,392,218,275,423,277,181,221,-200,-934,-933,-63,526,156,-502,-536,-7,306,52,-322,-398,-277,-89,127,70,-292,-253,443,817,258,-338,-235,-71,-424,-763,-596,-179,212,479,382,-22,-182,59,205,48,-116,-225,-359,-225,256,413,-99,-490,-118,381,266,-27,146,425,230,-216,-464,-497,-321,77,256,-62,-269,51,174,-362,-701,-294,-2,-435,-867,-679,-270,-11,251,492,435,94,-224,-303,-230,-300,-499,-421,-155,-292,-542,3,813,525,-378,-356,236,59,-440,-158,360,213,-159,-213,-224,-283,-187,-102,-26,397,852,617,-40,-251,59,325,245,-77,-271,-68,257,372,431,405,8,-215,399,931,275,-643,-517,98,254,134,-71,-397,-294,278,286,-310,-374,-9,-166,-455,-242,-196,-534,-388,67,-71,-327,12,279,131,288,559,151,-371,-259,-146,-390,-325,-80,-362,-695,-360,205,542,766,671,284,331,626,193,-439,-86,477,21,-594,-290,198,195,194,213,-202,-564,-309,1,-132,-285,-94,285,518,177,-638,-874,-54,667,393,-115,-67,173,196,122,-13,-165,-62,203,212,-6,-121,-109,-62,-20,-143,-350,-213,188,241,-56,-139,-30,-97,-103,249,531,395,244,337,230,-306,-715,-532,-147,-139,-283,70,753,841,134,-441,-250,245,427,308,153,103,215,343,235,23,72,257,174,-34,66,351,363,65,-263,-465,-462,-256,-32,133,278,113,-502,-738,8,605,-47,-727,25,1023,590,-277,42,744,454,-186,-132,141,17,-91,119,288,252,197,197,272,334,71,-455,-576,-92,275,50,-282,-159,219,278,-110,-464,-333,101,342,264,44,-171,-221,-31,135,92,134,411,451,-58,-643,-642,3,696,752,201,-169,11,161,-119,-356,-142,248,465,436,199,-35,-66,-114,-346,-377,-40,107,-149,-188,184,307,-18,-153,94,134,-159,-174,178,190,-319,-639,-448,-219,-213,-223,-179,-11,394,546,-4,-406,136,567,-95,-674,-118,536,461,336,272,-246,-483,247,783,319,-53,183,106,-249,31,576,509,151,5,-115,-94,288,421,-84,-479,-251,94,127,-22,-132,12,309,185,-329,-303,370,612,150,-129,25,61,-54,-11,49,-20,-28,34,4,-32,15,19,-25,-3,24,-12,-15,19,2,-19,9,12,-16,-2,16,-7,-11,13,2,-14,6,10,-11,-3,12,-5,-9,9,3,-11,4,8,-8,-3,9,-3,-7,7,3,-8,2,7,-6,-3,8,-1,-6,5,3,-7,1,6,-4,-3,6,0,-6,4,3,-5,0,5,-3,-3,5,0,-5,3,3,-4,-1,5,-2,-3,4,1,-4,2,3,-3,-1,4,-1,-3,3,1,-4,1,3,-3,-1,3,-1,-3,2,1,-3,0,3,-2,-2,3,0,-3,2,2,-2,0,2,-1,-2,2,0,-2,1,1,-2,0,2,-1,-1,2,0,-2,1,1,-1,-1,2,0,-1,1,1,-2,0,1,-1,-1,1,0,-1,1,1,-1,0,1,-1,-1,1,0,-1,1,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,1,0,-1,0,1,-1,0,1,0,-1,0,0,-1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- A saída da convolução vai ter tamanho 1572, mas só preciso dos 1060
	------------------------------------------------------------------------------

	-- TAMANHO 1572 - Símbolo OFDM parte real, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,-8,-252,-50,257,131,-90,5,157,127,28,-93,-149,13,112,-163,-382,-122,189,158,75,50,-166,-386,-280,-62,56,178,156,-138,-239,35,83,-201,-143,231,201,-134,-148,1,-117,-248,-126,-9,2,87,129,-59,-271,-297,-202,-33,141,83,-163,-215,-66,-97,-263,-163,123,159,-20,-31,131,200,217,341,368,100,-137,-28,131,38,-18,179,270,60,-114,-110,-115,-81,52,-8,-247,-187,132,176,39,121,92,-338,-512,-44,336,189,63,176,112,-90,-67,20,-13,69,172,-87,-376,-133,229,58,-304,-288,-133,-161,-152,-17,-24,-148,-149,-103,-160,-203,-158,-129,-90,43,175,221,202,51,-220,-289,-14,210,91,-72,3,85,-48,-167,-25,196,187,-7,-75,77,226,197,58,-77,-135,-26,191,227,19,-99,13,48,-119,-185,-14,138,105,-7,-104,-172,-151,2,184,210,29,-159,-169,-116,-120,-8,225,186,-104,-43,339,272,-225,-285,114,187,-14,158,477,337,16,45,179,45,-156,-171,-75,31,77,-34,-202,-229,-164,-112,-2,112,34,-119,-49,160,181,4,-106,-8,186,250,115,-8,-1,-61,-202,-102,179,155,-121,-81,239,290,115,159,267,41,-228,-63,287,284,-20,-204,-157,-101,-174,-232,-56,255,328,94,-53,36,11,-217,-228,49,140,-45,-60,109,12,-313,-394,-226,-153,-178,-138,-96,-73,16,11,-215,-365,-244,-130,-145,-76,-21,-204,-296,-6,207,-5,-209,-135,-115,-189,-86,-34,-244,-209,268,447,71,-90,178,183,-131,-134,82,-16,-223,-157,-133,-348,-375,-130,-45,-77,99,201,-86,-292,-7,338,313,117,-46,-220,-281,-96,99,58,-109,-215,-183,-6,125,-24,-241,-108,242,305,42,-131,-13,202,265,149,52,97,127,35,-9,56,57,36,179,300,140,-77,-95,-73,-87,46,211,125,-25,51,150,39,-51,65,170,68,-127,-204,-96,53,96,145,303,322,100,17,194,195,-36,-18,230,190,-114,-226,-86,105,261,236,-21,-195,-152,-181,-259,-17,368,361,41,-120,-67,-9,-6,-78,-192,-174,-20,54,55,143,232,174,56,-12,-31,-25,-94,-263,-259,57,301,220,109,115,43,-34,58,80,-61,3,278,314,123,46,8,-77,3,84,-165,-312,105,468,163,-240,-149,16,-107,-151,49,138,24,-13,76,92,-11,-104,-147,-217,-276,-153,82,98,-75,-58,66,-105,-355,-225,-21,-172,-298,-93,-26,-247,-185,209,309,60,-46,9,-52,-124,-38,49,49,107,235,277,184,49,-38,-69,-84,-63,5,-31,-274,-466,-325,-17,123,71,17,49,98,34,-101,-70,110,102,-80,-38,214,310,278,276,106,-174,-120,118,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- TAMANHO 1572 - Símbolo OFDM parte imaginária, -512 to 511
	--constant NOISY_ARRAY : T_NOISY_INPUT := (
	--	265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,-241,-142,-79,-110,-46,-71,-296,-384,-232,-109,17,300,443,217,-3,66,131,-16,-132,-64,31,78,150,181,59,-55,59,201,8,-327,-267,80,90,-225,-240,70,115,-147,-184,64,136,-73,-201,-68,116,121,0,-46,19,12,-155,-341,-401,-342,-250,-197,-172,-110,-78,-175,-203,51,280,108,-189,-172,11,80,137,199,80,-51,88,265,191,87,129,79,-124,-203,-104,-26,-33,-85,-129,-47,129,164,58,44,92,53,53,139,59,-177,-251,-176,-158,-81,88,14,-268,-254,66,195,108,138,211,138,91,111,-100,-466,-465,-32,262,78,-250,-268,-3,153,26,-161,-198,-138,-45,63,35,-146,-126,222,407,129,-168,-117,-36,-211,-380,-298,-89,106,239,191,-11,-91,29,102,24,-58,-112,-179,-112,128,206,-49,-245,-59,190,133,-14,73,212,114,-108,-231,-248,-160,38,128,-31,-134,26,87,-180,-350,-147,-1,-217,-432,-339,-134,-5,125,246,217,47,-112,-151,-115,-150,-249,-210,-77,-146,-270,1,405,262,-189,-178,118,30,-220,-79,180,106,-79,-106,-112,-141,-93,-51,-13,198,425,308,-20,-125,29,162,122,-38,-135,-34,128,186,215,202,4,-107,199,465,137,-321,-258,49,127,67,-36,-198,-147,139,143,-155,-187,-4,-83,-227,-121,-98,-266,-193,34,-35,-163,6,139,66,144,279,76,-185,-129,-73,-194,-162,-40,-181,-347,-180,102,270,382,335,142,165,312,96,-219,-43,238,11,-296,-145,99,97,97,106,-101,-281,-154,1,-66,-142,-47,142,258,89,-318,-436,-27,333,196,-58,-33,86,98,61,-7,-83,-31,102,105,-3,-60,-55,-31,-10,-72,-175,-106,94,120,-28,-69,-15,-49,-51,124,265,197,122,168,114,-152,-357,-266,-73,-69,-142,35,376,419,67,-220,-125,122,213,154,76,51,108,171,117,12,36,128,87,-17,32,175,182,32,-132,-231,-230,-128,-16,67,138,56,-250,-368,3,302,-23,-363,13,511,294,-139,22,371,226,-92,-65,70,9,-45,59,143,127,98,97,136,167,34,-227,-286,-46,137,26,-140,-81,110,140,-56,-232,-165,50,170,133,23,-87,-110,-14,66,45,69,205,223,-28,-320,-322,2,349,374,100,-83,5,79,-58,-176,-73,124,234,216,98,-15,-33,-59,-171,-187,-22,53,-71,-95,90,156,-9,-79,48,69,-82,-88,92,94,-162,-316,-222,-113,-105,-108,-92,-7,200,271,-5,-199,70,278,-47,-332,-62,265,235,167,131,-119,-238,118,391,165,-30,88,59,-124,9,292,259,68,2,-49,-52,137,219,-41,-250,-120,55,52,-13,-50,-1,141,111,-159,-179,199,340,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0	
	--);
	-- A saída da convolução vai ter tamanho 2596, mas só preciso dos 1572
	
	component fir_filter_lms
	port (
		clk      : in  std_logic   ;
		reset    : in  std_logic   ;
		i_data   : in  IN_TYPE	   ;
		i_ref    : in  IN_TYPE	   ;
		o_coeff1 : out IN_TYPE     ;
		o_coeff2 : out IN_TYPE     ;
		o_data   : out OUT_TYPE    ;
		o_error  : out OUT_TYPE    );
	end component;

	signal i_data   : IN_TYPE;
	signal i_ref   : IN_TYPE;
	signal NOISY	: ARRAY_COEFF(0 to noisy_size-1);
	signal NOISYF	: ARRAY_COEFF(0 to noisy_size-1);

begin
	
	u_fir_filter_lms : fir_filter_lms
	port map(
		clk         => clk       	,
		reset       => reset      	,
		i_data      => i_data 		,
		i_ref       => i_ref 		,
		o_coeff1     => o_fir_coeff1 		,
		o_coeff2     => o_fir_coeff2 		,
		o_data     	=> o_data_buffer ,
		o_error     => o_error       );

	p_input : process (reset,clk)
		variable control  	: unsigned(11 downto 0):= (others=>'0');
		variable count 		: integer := 0;
		variable count2     : integer := 0;
		variable s			: integer RANGE 0 TO 2**8-1 :=255;
		variable first_time : std_logic := '0';
	begin
		if(reset=BUTTON_HIGH) then
			i_data      <= (others=>'0'); 
			i_ref       <= (others=>'0'); 
			count 		:= 0;
			count2 		:= 0;
			first_time	:='0';
		elsif(falling_edge(clk)) then
			if(first_time='0') then
				for k in 0 to noisy_size-1 loop
					NOISYF(k)  <=  std_logic_vector(to_signed(NOISYF_ARRAY(k),Win));
				end loop;			
				for j in 0 to noisy_size-1 loop
					NOISY(j)  <=  std_logic_vector(to_signed(NOISY_ARRAY(j),Win));
				end loop;
				first_time := '1';
			else
				
				-- NOISY ANALOG SIGNAL
				if(count < noisy_size) then
					i_data <= NOISY(count);
					i_ref <= NOISYF(count);					
					count := count + 1;
				else
					i_data <= (others=>'0');
					i_ref <= (others=>'0');
				end if;
				-------------------------------------------------

				-- COEFFICIENTS
				--if(count < Lfilter-1) then
				--	o_fir_coeff <= o_coeff(count);
				--else
				--	o_fir_coeff <= (others=>'0');
				--end if;
				---------------------------------------------------
				o_inputref <= i_ref;
				o_inputdata <= i_data;
				--count := count+1;
			end if;
		end if;
	end process p_input;





end rtl;
